module cc_dir_ext( // @[:anonymous source@2.2]
  input  [9:0]   RW0_addr, // @[:anonymous source@3.4]
  input          RW0_clk, // @[:anonymous source@4.4]
  input  [127:0] RW0_wdata, // @[:anonymous source@5.4]
  output [127:0] RW0_rdata, // @[:anonymous source@6.4]
  input          RW0_en, // @[:anonymous source@7.4]
  input          RW0_wmode, // @[:anonymous source@8.4]
  input  [7:0]   RW0_wmask // @[:anonymous source@9.4]
);
  wire [9:0] mem_0_0_RW0_addr; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@11.4]
  wire [15:0] mem_0_0_RW0_wdata; // @[:anonymous source@11.4]
  wire [15:0] mem_0_0_RW0_rdata; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@11.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@11.4]
  wire [9:0] mem_0_1_RW0_addr; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@12.4]
  wire [15:0] mem_0_1_RW0_wdata; // @[:anonymous source@12.4]
  wire [15:0] mem_0_1_RW0_rdata; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@12.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@12.4]
  wire [9:0] mem_0_2_RW0_addr; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@13.4]
  wire [15:0] mem_0_2_RW0_wdata; // @[:anonymous source@13.4]
  wire [15:0] mem_0_2_RW0_rdata; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@13.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@13.4]
  wire [9:0] mem_0_3_RW0_addr; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@14.4]
  wire [15:0] mem_0_3_RW0_wdata; // @[:anonymous source@14.4]
  wire [15:0] mem_0_3_RW0_rdata; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@14.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@14.4]
  wire [9:0] mem_0_4_RW0_addr; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_clk; // @[:anonymous source@15.4]
  wire [15:0] mem_0_4_RW0_wdata; // @[:anonymous source@15.4]
  wire [15:0] mem_0_4_RW0_rdata; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_en; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_wmode; // @[:anonymous source@15.4]
  wire  mem_0_4_RW0_wmask; // @[:anonymous source@15.4]
  wire [9:0] mem_0_5_RW0_addr; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_clk; // @[:anonymous source@16.4]
  wire [15:0] mem_0_5_RW0_wdata; // @[:anonymous source@16.4]
  wire [15:0] mem_0_5_RW0_rdata; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_en; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_wmode; // @[:anonymous source@16.4]
  wire  mem_0_5_RW0_wmask; // @[:anonymous source@16.4]
  wire [9:0] mem_0_6_RW0_addr; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_clk; // @[:anonymous source@17.4]
  wire [15:0] mem_0_6_RW0_wdata; // @[:anonymous source@17.4]
  wire [15:0] mem_0_6_RW0_rdata; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_en; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_wmode; // @[:anonymous source@17.4]
  wire  mem_0_6_RW0_wmask; // @[:anonymous source@17.4]
  wire [9:0] mem_0_7_RW0_addr; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_clk; // @[:anonymous source@18.4]
  wire [15:0] mem_0_7_RW0_wdata; // @[:anonymous source@18.4]
  wire [15:0] mem_0_7_RW0_rdata; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_en; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_wmode; // @[:anonymous source@18.4]
  wire  mem_0_7_RW0_wmask; // @[:anonymous source@18.4]
  wire [15:0] RW0_rdata_0_0; // @[:anonymous source@21.4]
  wire [15:0] RW0_rdata_0_1; // @[:anonymous source@28.4]
  wire [15:0] RW0_rdata_0_2; // @[:anonymous source@35.4]
  wire [15:0] RW0_rdata_0_3; // @[:anonymous source@42.4]
  wire [15:0] RW0_rdata_0_4; // @[:anonymous source@49.4]
  wire [15:0] RW0_rdata_0_5; // @[:anonymous source@56.4]
  wire [15:0] RW0_rdata_0_6; // @[:anonymous source@63.4]
  wire [15:0] RW0_rdata_0_7; // @[:anonymous source@70.4]
  wire [31:0] _GEN_0; // @[:anonymous source@75.4]
  wire [47:0] _GEN_1; // @[:anonymous source@75.4]
  wire [63:0] _GEN_2; // @[:anonymous source@75.4]
  wire [79:0] _GEN_3; // @[:anonymous source@75.4]
  wire [95:0] _GEN_4; // @[:anonymous source@75.4]
  wire [111:0] _GEN_5; // @[:anonymous source@75.4]
  wire [127:0] RW0_rdata_0; // @[:anonymous source@75.4]
  wire [31:0] _GEN_6; // @[:anonymous source@76.4]
  wire [47:0] _GEN_7; // @[:anonymous source@76.4]
  wire [63:0] _GEN_8; // @[:anonymous source@76.4]
  wire [79:0] _GEN_9; // @[:anonymous source@76.4]
  wire [95:0] _GEN_10; // @[:anonymous source@76.4]
  wire [111:0] _GEN_11; // @[:anonymous source@76.4]
  split_cc_dir_ext mem_0_0 ( // @[:anonymous source@11.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_cc_dir_ext mem_0_1 ( // @[:anonymous source@12.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_cc_dir_ext mem_0_2 ( // @[:anonymous source@13.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_cc_dir_ext mem_0_3 ( // @[:anonymous source@14.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  split_cc_dir_ext mem_0_4 ( // @[:anonymous source@15.4]
    .RW0_addr(mem_0_4_RW0_addr),
    .RW0_clk(mem_0_4_RW0_clk),
    .RW0_wdata(mem_0_4_RW0_wdata),
    .RW0_rdata(mem_0_4_RW0_rdata),
    .RW0_en(mem_0_4_RW0_en),
    .RW0_wmode(mem_0_4_RW0_wmode),
    .RW0_wmask(mem_0_4_RW0_wmask)
  );
  split_cc_dir_ext mem_0_5 ( // @[:anonymous source@16.4]
    .RW0_addr(mem_0_5_RW0_addr),
    .RW0_clk(mem_0_5_RW0_clk),
    .RW0_wdata(mem_0_5_RW0_wdata),
    .RW0_rdata(mem_0_5_RW0_rdata),
    .RW0_en(mem_0_5_RW0_en),
    .RW0_wmode(mem_0_5_RW0_wmode),
    .RW0_wmask(mem_0_5_RW0_wmask)
  );
  split_cc_dir_ext mem_0_6 ( // @[:anonymous source@17.4]
    .RW0_addr(mem_0_6_RW0_addr),
    .RW0_clk(mem_0_6_RW0_clk),
    .RW0_wdata(mem_0_6_RW0_wdata),
    .RW0_rdata(mem_0_6_RW0_rdata),
    .RW0_en(mem_0_6_RW0_en),
    .RW0_wmode(mem_0_6_RW0_wmode),
    .RW0_wmask(mem_0_6_RW0_wmask)
  );
  split_cc_dir_ext mem_0_7 ( // @[:anonymous source@18.4]
    .RW0_addr(mem_0_7_RW0_addr),
    .RW0_clk(mem_0_7_RW0_clk),
    .RW0_wdata(mem_0_7_RW0_wdata),
    .RW0_rdata(mem_0_7_RW0_rdata),
    .RW0_en(mem_0_7_RW0_en),
    .RW0_wmode(mem_0_7_RW0_wmode),
    .RW0_wmask(mem_0_7_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@21.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@28.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@35.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@42.4]
  assign RW0_rdata_0_4 = mem_0_4_RW0_rdata; // @[:anonymous source@49.4]
  assign RW0_rdata_0_5 = mem_0_5_RW0_rdata; // @[:anonymous source@56.4]
  assign RW0_rdata_0_6 = mem_0_6_RW0_rdata; // @[:anonymous source@63.4]
  assign RW0_rdata_0_7 = mem_0_7_RW0_rdata; // @[:anonymous source@70.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_2 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_3 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_4 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_5 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign RW0_rdata_0 = {RW0_rdata_0_7,RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@75.4]
  assign _GEN_6 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_7 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_8 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_9 = {RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_10 = {RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign _GEN_11 = {RW0_rdata_0_6,RW0_rdata_0_5,RW0_rdata_0_4,RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@76.4]
  assign RW0_rdata = {RW0_rdata_0_7,_GEN_5}; // @[:anonymous source@76.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@20.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@19.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[15:0]; // @[:anonymous source@22.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@25.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@24.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@23.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@27.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@26.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[31:16]; // @[:anonymous source@29.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@32.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@31.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@30.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@34.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@33.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[47:32]; // @[:anonymous source@36.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@39.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@38.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@37.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@41.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@40.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[63:48]; // @[:anonymous source@43.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@46.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@45.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@44.4]
  assign mem_0_4_RW0_addr = RW0_addr; // @[:anonymous source@48.4]
  assign mem_0_4_RW0_clk = RW0_clk; // @[:anonymous source@47.4]
  assign mem_0_4_RW0_wdata = RW0_wdata[79:64]; // @[:anonymous source@50.4]
  assign mem_0_4_RW0_en = RW0_en; // @[:anonymous source@53.4]
  assign mem_0_4_RW0_wmode = RW0_wmode; // @[:anonymous source@52.4]
  assign mem_0_4_RW0_wmask = RW0_wmask[4]; // @[:anonymous source@51.4]
  assign mem_0_5_RW0_addr = RW0_addr; // @[:anonymous source@55.4]
  assign mem_0_5_RW0_clk = RW0_clk; // @[:anonymous source@54.4]
  assign mem_0_5_RW0_wdata = RW0_wdata[95:80]; // @[:anonymous source@57.4]
  assign mem_0_5_RW0_en = RW0_en; // @[:anonymous source@60.4]
  assign mem_0_5_RW0_wmode = RW0_wmode; // @[:anonymous source@59.4]
  assign mem_0_5_RW0_wmask = RW0_wmask[5]; // @[:anonymous source@58.4]
  assign mem_0_6_RW0_addr = RW0_addr; // @[:anonymous source@62.4]
  assign mem_0_6_RW0_clk = RW0_clk; // @[:anonymous source@61.4]
  assign mem_0_6_RW0_wdata = RW0_wdata[111:96]; // @[:anonymous source@64.4]
  assign mem_0_6_RW0_en = RW0_en; // @[:anonymous source@67.4]
  assign mem_0_6_RW0_wmode = RW0_wmode; // @[:anonymous source@66.4]
  assign mem_0_6_RW0_wmask = RW0_wmask[6]; // @[:anonymous source@65.4]
  assign mem_0_7_RW0_addr = RW0_addr; // @[:anonymous source@69.4]
  assign mem_0_7_RW0_clk = RW0_clk; // @[:anonymous source@68.4]
  assign mem_0_7_RW0_wdata = RW0_wdata[127:112]; // @[:anonymous source@71.4]
  assign mem_0_7_RW0_en = RW0_en; // @[:anonymous source@74.4]
  assign mem_0_7_RW0_wmode = RW0_wmode; // @[:anonymous source@73.4]
  assign mem_0_7_RW0_wmask = RW0_wmask[7]; // @[:anonymous source@72.4]
endmodule
module cc_banks_0_ext( // @[:anonymous source@78.2]
  input  [13:0] RW0_addr, // @[:anonymous source@79.4]
  input         RW0_clk, // @[:anonymous source@80.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@81.4]
  output [63:0] RW0_rdata, // @[:anonymous source@82.4]
  input         RW0_en, // @[:anonymous source@83.4]
  input         RW0_wmode // @[:anonymous source@84.4]
);
  wire [13:0] mem_0_0_RW0_addr; // @[:anonymous source@86.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@86.4]
  wire [63:0] mem_0_0_RW0_wdata; // @[:anonymous source@86.4]
  wire [63:0] mem_0_0_RW0_rdata; // @[:anonymous source@86.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@86.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@86.4]
  wire [63:0] RW0_rdata_0_0; // @[:anonymous source@89.4]
  wire [63:0] RW0_rdata_0; // @[:anonymous source@93.4]
  split_cc_banks_0_ext mem_0_0 ( // @[:anonymous source@86.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@89.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@93.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@94.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@88.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@87.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@90.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@92.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@91.4]
endmodule
module tag_array_ext( // @[:anonymous source@96.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@97.4]
  input         RW0_clk, // @[:anonymous source@98.4]
  input  [87:0] RW0_wdata, // @[:anonymous source@99.4]
  output [87:0] RW0_rdata, // @[:anonymous source@100.4]
  input         RW0_en, // @[:anonymous source@101.4]
  input         RW0_wmode, // @[:anonymous source@102.4]
  input  [3:0]  RW0_wmask // @[:anonymous source@103.4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@105.4]
  wire [21:0] mem_0_0_RW0_wdata; // @[:anonymous source@105.4]
  wire [21:0] mem_0_0_RW0_rdata; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@105.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@105.4]
  wire [5:0] mem_0_1_RW0_addr; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@106.4]
  wire [21:0] mem_0_1_RW0_wdata; // @[:anonymous source@106.4]
  wire [21:0] mem_0_1_RW0_rdata; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@106.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@106.4]
  wire [5:0] mem_0_2_RW0_addr; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@107.4]
  wire [21:0] mem_0_2_RW0_wdata; // @[:anonymous source@107.4]
  wire [21:0] mem_0_2_RW0_rdata; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@107.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@107.4]
  wire [5:0] mem_0_3_RW0_addr; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@108.4]
  wire [21:0] mem_0_3_RW0_wdata; // @[:anonymous source@108.4]
  wire [21:0] mem_0_3_RW0_rdata; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@108.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@108.4]
  wire [21:0] RW0_rdata_0_0; // @[:anonymous source@111.4]
  wire [21:0] RW0_rdata_0_1; // @[:anonymous source@118.4]
  wire [21:0] RW0_rdata_0_2; // @[:anonymous source@125.4]
  wire [21:0] RW0_rdata_0_3; // @[:anonymous source@132.4]
  wire [43:0] _GEN_0; // @[:anonymous source@137.4]
  wire [65:0] _GEN_1; // @[:anonymous source@137.4]
  wire [87:0] RW0_rdata_0; // @[:anonymous source@137.4]
  wire [43:0] _GEN_2; // @[:anonymous source@138.4]
  wire [65:0] _GEN_3; // @[:anonymous source@138.4]
  split_tag_array_ext mem_0_0 ( // @[:anonymous source@105.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_ext mem_0_1 ( // @[:anonymous source@106.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_ext mem_0_2 ( // @[:anonymous source@107.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_ext mem_0_3 ( // @[:anonymous source@108.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@111.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@118.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@125.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@132.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@137.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@137.4]
  assign RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@137.4]
  assign _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@138.4]
  assign _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@138.4]
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[:anonymous source@138.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@110.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@109.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[21:0]; // @[:anonymous source@112.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@115.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@114.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@113.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@117.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@116.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[43:22]; // @[:anonymous source@119.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@122.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@121.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@120.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@124.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@123.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[65:44]; // @[:anonymous source@126.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@129.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@128.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@127.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@131.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@130.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[87:66]; // @[:anonymous source@133.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@136.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@135.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@134.4]
endmodule
module array_0_0_ext( // @[:anonymous source@140.2]
  input  [8:0]  W0_addr, // @[:anonymous source@141.4]
  input         W0_clk, // @[:anonymous source@142.4]
  input  [63:0] W0_data, // @[:anonymous source@143.4]
  input         W0_en, // @[:anonymous source@144.4]
  input         W0_mask, // @[:anonymous source@145.4]
  input  [8:0]  R0_addr, // @[:anonymous source@146.4]
  input         R0_clk, // @[:anonymous source@147.4]
  output [63:0] R0_data, // @[:anonymous source@148.4]
  input         R0_en // @[:anonymous source@149.4]
);
  wire [8:0] mem_0_0_W0_addr; // @[:anonymous source@151.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@151.4]
  wire [63:0] mem_0_0_W0_data; // @[:anonymous source@151.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@151.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@151.4]
  wire [8:0] mem_0_0_R0_addr; // @[:anonymous source@151.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@151.4]
  wire [63:0] mem_0_0_R0_data; // @[:anonymous source@151.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@151.4]
  wire [63:0] R0_data_0_0; // @[:anonymous source@159.4]
  wire [63:0] R0_data_0; // @[:anonymous source@161.4]
  split_array_0_0_ext mem_0_0 ( // @[:anonymous source@151.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@159.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@161.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@162.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@153.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@152.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@154.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@156.4]
  assign mem_0_0_W0_mask = W0_mask; // @[:anonymous source@155.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@158.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@157.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@160.4]
endmodule
module tag_array_0_ext( // @[:anonymous source@164.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@165.4]
  input         RW0_clk, // @[:anonymous source@166.4]
  input  [79:0] RW0_wdata, // @[:anonymous source@167.4]
  output [79:0] RW0_rdata, // @[:anonymous source@168.4]
  input         RW0_en, // @[:anonymous source@169.4]
  input         RW0_wmode, // @[:anonymous source@170.4]
  input  [3:0]  RW0_wmask // @[:anonymous source@171.4]
);
  wire [5:0] mem_0_0_RW0_addr; // @[:anonymous source@173.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@173.4]
  wire [19:0] mem_0_0_RW0_wdata; // @[:anonymous source@173.4]
  wire [19:0] mem_0_0_RW0_rdata; // @[:anonymous source@173.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@173.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@173.4]
  wire  mem_0_0_RW0_wmask; // @[:anonymous source@173.4]
  wire [5:0] mem_0_1_RW0_addr; // @[:anonymous source@174.4]
  wire  mem_0_1_RW0_clk; // @[:anonymous source@174.4]
  wire [19:0] mem_0_1_RW0_wdata; // @[:anonymous source@174.4]
  wire [19:0] mem_0_1_RW0_rdata; // @[:anonymous source@174.4]
  wire  mem_0_1_RW0_en; // @[:anonymous source@174.4]
  wire  mem_0_1_RW0_wmode; // @[:anonymous source@174.4]
  wire  mem_0_1_RW0_wmask; // @[:anonymous source@174.4]
  wire [5:0] mem_0_2_RW0_addr; // @[:anonymous source@175.4]
  wire  mem_0_2_RW0_clk; // @[:anonymous source@175.4]
  wire [19:0] mem_0_2_RW0_wdata; // @[:anonymous source@175.4]
  wire [19:0] mem_0_2_RW0_rdata; // @[:anonymous source@175.4]
  wire  mem_0_2_RW0_en; // @[:anonymous source@175.4]
  wire  mem_0_2_RW0_wmode; // @[:anonymous source@175.4]
  wire  mem_0_2_RW0_wmask; // @[:anonymous source@175.4]
  wire [5:0] mem_0_3_RW0_addr; // @[:anonymous source@176.4]
  wire  mem_0_3_RW0_clk; // @[:anonymous source@176.4]
  wire [19:0] mem_0_3_RW0_wdata; // @[:anonymous source@176.4]
  wire [19:0] mem_0_3_RW0_rdata; // @[:anonymous source@176.4]
  wire  mem_0_3_RW0_en; // @[:anonymous source@176.4]
  wire  mem_0_3_RW0_wmode; // @[:anonymous source@176.4]
  wire  mem_0_3_RW0_wmask; // @[:anonymous source@176.4]
  wire [19:0] RW0_rdata_0_0; // @[:anonymous source@179.4]
  wire [19:0] RW0_rdata_0_1; // @[:anonymous source@186.4]
  wire [19:0] RW0_rdata_0_2; // @[:anonymous source@193.4]
  wire [19:0] RW0_rdata_0_3; // @[:anonymous source@200.4]
  wire [39:0] _GEN_0; // @[:anonymous source@205.4]
  wire [59:0] _GEN_1; // @[:anonymous source@205.4]
  wire [79:0] RW0_rdata_0; // @[:anonymous source@205.4]
  wire [39:0] _GEN_2; // @[:anonymous source@206.4]
  wire [59:0] _GEN_3; // @[:anonymous source@206.4]
  split_tag_array_0_ext mem_0_0 ( // @[:anonymous source@173.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_1 ( // @[:anonymous source@174.4]
    .RW0_addr(mem_0_1_RW0_addr),
    .RW0_clk(mem_0_1_RW0_clk),
    .RW0_wdata(mem_0_1_RW0_wdata),
    .RW0_rdata(mem_0_1_RW0_rdata),
    .RW0_en(mem_0_1_RW0_en),
    .RW0_wmode(mem_0_1_RW0_wmode),
    .RW0_wmask(mem_0_1_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_2 ( // @[:anonymous source@175.4]
    .RW0_addr(mem_0_2_RW0_addr),
    .RW0_clk(mem_0_2_RW0_clk),
    .RW0_wdata(mem_0_2_RW0_wdata),
    .RW0_rdata(mem_0_2_RW0_rdata),
    .RW0_en(mem_0_2_RW0_en),
    .RW0_wmode(mem_0_2_RW0_wmode),
    .RW0_wmask(mem_0_2_RW0_wmask)
  );
  split_tag_array_0_ext mem_0_3 ( // @[:anonymous source@176.4]
    .RW0_addr(mem_0_3_RW0_addr),
    .RW0_clk(mem_0_3_RW0_clk),
    .RW0_wdata(mem_0_3_RW0_wdata),
    .RW0_rdata(mem_0_3_RW0_rdata),
    .RW0_en(mem_0_3_RW0_en),
    .RW0_wmode(mem_0_3_RW0_wmode),
    .RW0_wmask(mem_0_3_RW0_wmask)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@179.4]
  assign RW0_rdata_0_1 = mem_0_1_RW0_rdata; // @[:anonymous source@186.4]
  assign RW0_rdata_0_2 = mem_0_2_RW0_rdata; // @[:anonymous source@193.4]
  assign RW0_rdata_0_3 = mem_0_3_RW0_rdata; // @[:anonymous source@200.4]
  assign _GEN_0 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@205.4]
  assign _GEN_1 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@205.4]
  assign RW0_rdata_0 = {RW0_rdata_0_3,RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@205.4]
  assign _GEN_2 = {RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@206.4]
  assign _GEN_3 = {RW0_rdata_0_2,RW0_rdata_0_1,RW0_rdata_0_0}; // @[:anonymous source@206.4]
  assign RW0_rdata = {RW0_rdata_0_3,_GEN_1}; // @[:anonymous source@206.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@178.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@177.4]
  assign mem_0_0_RW0_wdata = RW0_wdata[19:0]; // @[:anonymous source@180.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@183.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@182.4]
  assign mem_0_0_RW0_wmask = RW0_wmask[0]; // @[:anonymous source@181.4]
  assign mem_0_1_RW0_addr = RW0_addr; // @[:anonymous source@185.4]
  assign mem_0_1_RW0_clk = RW0_clk; // @[:anonymous source@184.4]
  assign mem_0_1_RW0_wdata = RW0_wdata[39:20]; // @[:anonymous source@187.4]
  assign mem_0_1_RW0_en = RW0_en; // @[:anonymous source@190.4]
  assign mem_0_1_RW0_wmode = RW0_wmode; // @[:anonymous source@189.4]
  assign mem_0_1_RW0_wmask = RW0_wmask[1]; // @[:anonymous source@188.4]
  assign mem_0_2_RW0_addr = RW0_addr; // @[:anonymous source@192.4]
  assign mem_0_2_RW0_clk = RW0_clk; // @[:anonymous source@191.4]
  assign mem_0_2_RW0_wdata = RW0_wdata[59:40]; // @[:anonymous source@194.4]
  assign mem_0_2_RW0_en = RW0_en; // @[:anonymous source@197.4]
  assign mem_0_2_RW0_wmode = RW0_wmode; // @[:anonymous source@196.4]
  assign mem_0_2_RW0_wmask = RW0_wmask[2]; // @[:anonymous source@195.4]
  assign mem_0_3_RW0_addr = RW0_addr; // @[:anonymous source@199.4]
  assign mem_0_3_RW0_clk = RW0_clk; // @[:anonymous source@198.4]
  assign mem_0_3_RW0_wdata = RW0_wdata[79:60]; // @[:anonymous source@201.4]
  assign mem_0_3_RW0_en = RW0_en; // @[:anonymous source@204.4]
  assign mem_0_3_RW0_wmode = RW0_wmode; // @[:anonymous source@203.4]
  assign mem_0_3_RW0_wmask = RW0_wmask[3]; // @[:anonymous source@202.4]
endmodule
module dataArrayWay_0_ext( // @[:anonymous source@208.2]
  input  [8:0]  RW0_addr, // @[:anonymous source@209.4]
  input         RW0_clk, // @[:anonymous source@210.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@211.4]
  output [63:0] RW0_rdata, // @[:anonymous source@212.4]
  input         RW0_en, // @[:anonymous source@213.4]
  input         RW0_wmode // @[:anonymous source@214.4]
);
  wire [8:0] mem_0_0_RW0_addr; // @[:anonymous source@216.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@216.4]
  wire [63:0] mem_0_0_RW0_wdata; // @[:anonymous source@216.4]
  wire [63:0] mem_0_0_RW0_rdata; // @[:anonymous source@216.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@216.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@216.4]
  wire [63:0] RW0_rdata_0_0; // @[:anonymous source@219.4]
  wire [63:0] RW0_rdata_0; // @[:anonymous source@223.4]
  split_dataArrayWay_0_ext mem_0_0 ( // @[:anonymous source@216.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@219.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@223.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@224.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@218.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@217.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@220.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@222.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@221.4]
endmodule
module hi_us_ext( // @[:anonymous source@226.2]
  input  [6:0] W0_addr, // @[:anonymous source@227.4]
  input        W0_clk, // @[:anonymous source@228.4]
  input  [3:0] W0_data, // @[:anonymous source@229.4]
  input        W0_en, // @[:anonymous source@230.4]
  input  [3:0] W0_mask, // @[:anonymous source@231.4]
  input  [6:0] R0_addr, // @[:anonymous source@232.4]
  input        R0_clk, // @[:anonymous source@233.4]
  output [3:0] R0_data, // @[:anonymous source@234.4]
  input        R0_en // @[:anonymous source@235.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@237.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@237.4]
  wire  mem_0_0_W0_data; // @[:anonymous source@237.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@237.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@237.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@237.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@237.4]
  wire  mem_0_0_R0_data; // @[:anonymous source@237.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@237.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@238.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@238.4]
  wire  mem_0_1_W0_data; // @[:anonymous source@238.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@238.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@238.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@238.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@238.4]
  wire  mem_0_1_R0_data; // @[:anonymous source@238.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@238.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@239.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@239.4]
  wire  mem_0_2_W0_data; // @[:anonymous source@239.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@239.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@239.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@239.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@239.4]
  wire  mem_0_2_R0_data; // @[:anonymous source@239.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@239.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@240.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@240.4]
  wire  mem_0_3_W0_data; // @[:anonymous source@240.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@240.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@240.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@240.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@240.4]
  wire  mem_0_3_R0_data; // @[:anonymous source@240.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@240.4]
  wire  R0_data_0_0; // @[:anonymous source@263.4]
  wire  R0_data_0_1; // @[:anonymous source@267.4]
  wire  R0_data_0_2; // @[:anonymous source@271.4]
  wire  R0_data_0_3; // @[:anonymous source@275.4]
  wire [1:0] _GEN_0; // @[:anonymous source@277.4]
  wire [2:0] _GEN_1; // @[:anonymous source@277.4]
  wire [3:0] R0_data_0; // @[:anonymous source@277.4]
  wire [1:0] _GEN_2; // @[:anonymous source@278.4]
  wire [2:0] _GEN_3; // @[:anonymous source@278.4]
  split_hi_us_ext mem_0_0 ( // @[:anonymous source@237.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_hi_us_ext mem_0_1 ( // @[:anonymous source@238.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_hi_us_ext mem_0_2 ( // @[:anonymous source@239.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_hi_us_ext mem_0_3 ( // @[:anonymous source@240.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@263.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@267.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@271.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@275.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@277.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@277.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@277.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@278.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@278.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@278.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@242.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@241.4]
  assign mem_0_0_W0_data = W0_data[0]; // @[:anonymous source@243.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@245.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@244.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@262.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@261.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@264.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@247.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@246.4]
  assign mem_0_1_W0_data = W0_data[1]; // @[:anonymous source@248.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@250.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@249.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@266.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@265.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@268.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@252.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@251.4]
  assign mem_0_2_W0_data = W0_data[2]; // @[:anonymous source@253.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@255.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@254.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@270.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@269.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@272.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@257.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@256.4]
  assign mem_0_3_W0_data = W0_data[3]; // @[:anonymous source@258.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@260.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@259.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@274.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@273.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@276.4]
endmodule
module table_ext( // @[:anonymous source@280.2]
  input  [6:0]  W0_addr, // @[:anonymous source@281.4]
  input         W0_clk, // @[:anonymous source@282.4]
  input  [43:0] W0_data, // @[:anonymous source@283.4]
  input         W0_en, // @[:anonymous source@284.4]
  input  [3:0]  W0_mask, // @[:anonymous source@285.4]
  input  [6:0]  R0_addr, // @[:anonymous source@286.4]
  input         R0_clk, // @[:anonymous source@287.4]
  output [43:0] R0_data, // @[:anonymous source@288.4]
  input         R0_en // @[:anonymous source@289.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@291.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@291.4]
  wire [10:0] mem_0_0_W0_data; // @[:anonymous source@291.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@291.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@291.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@291.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@291.4]
  wire [10:0] mem_0_0_R0_data; // @[:anonymous source@291.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@291.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@292.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@292.4]
  wire [10:0] mem_0_1_W0_data; // @[:anonymous source@292.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@292.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@292.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@292.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@292.4]
  wire [10:0] mem_0_1_R0_data; // @[:anonymous source@292.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@292.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@293.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@293.4]
  wire [10:0] mem_0_2_W0_data; // @[:anonymous source@293.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@293.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@293.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@293.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@293.4]
  wire [10:0] mem_0_2_R0_data; // @[:anonymous source@293.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@293.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@294.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@294.4]
  wire [10:0] mem_0_3_W0_data; // @[:anonymous source@294.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@294.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@294.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@294.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@294.4]
  wire [10:0] mem_0_3_R0_data; // @[:anonymous source@294.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@294.4]
  wire [10:0] R0_data_0_0; // @[:anonymous source@317.4]
  wire [10:0] R0_data_0_1; // @[:anonymous source@321.4]
  wire [10:0] R0_data_0_2; // @[:anonymous source@325.4]
  wire [10:0] R0_data_0_3; // @[:anonymous source@329.4]
  wire [21:0] _GEN_0; // @[:anonymous source@331.4]
  wire [32:0] _GEN_1; // @[:anonymous source@331.4]
  wire [43:0] R0_data_0; // @[:anonymous source@331.4]
  wire [21:0] _GEN_2; // @[:anonymous source@332.4]
  wire [32:0] _GEN_3; // @[:anonymous source@332.4]
  split_table_ext mem_0_0 ( // @[:anonymous source@291.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_table_ext mem_0_1 ( // @[:anonymous source@292.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_table_ext mem_0_2 ( // @[:anonymous source@293.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_table_ext mem_0_3 ( // @[:anonymous source@294.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@317.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@321.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@325.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@329.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@331.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@331.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@331.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@332.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@332.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@332.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@296.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@295.4]
  assign mem_0_0_W0_data = W0_data[10:0]; // @[:anonymous source@297.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@299.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@298.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@316.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@315.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@318.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@301.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@300.4]
  assign mem_0_1_W0_data = W0_data[21:11]; // @[:anonymous source@302.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@304.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@303.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@320.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@319.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@322.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@306.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@305.4]
  assign mem_0_2_W0_data = W0_data[32:22]; // @[:anonymous source@307.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@309.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@308.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@324.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@323.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@326.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@311.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@310.4]
  assign mem_0_3_W0_data = W0_data[43:33]; // @[:anonymous source@312.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@314.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@313.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@328.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@327.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@330.4]
endmodule
module hi_us_0_ext( // @[:anonymous source@334.2]
  input  [7:0] W0_addr, // @[:anonymous source@335.4]
  input        W0_clk, // @[:anonymous source@336.4]
  input  [3:0] W0_data, // @[:anonymous source@337.4]
  input        W0_en, // @[:anonymous source@338.4]
  input  [3:0] W0_mask, // @[:anonymous source@339.4]
  input  [7:0] R0_addr, // @[:anonymous source@340.4]
  input        R0_clk, // @[:anonymous source@341.4]
  output [3:0] R0_data, // @[:anonymous source@342.4]
  input        R0_en // @[:anonymous source@343.4]
);
  wire [7:0] mem_0_0_W0_addr; // @[:anonymous source@345.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@345.4]
  wire  mem_0_0_W0_data; // @[:anonymous source@345.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@345.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@345.4]
  wire [7:0] mem_0_0_R0_addr; // @[:anonymous source@345.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@345.4]
  wire  mem_0_0_R0_data; // @[:anonymous source@345.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@345.4]
  wire [7:0] mem_0_1_W0_addr; // @[:anonymous source@346.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@346.4]
  wire  mem_0_1_W0_data; // @[:anonymous source@346.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@346.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@346.4]
  wire [7:0] mem_0_1_R0_addr; // @[:anonymous source@346.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@346.4]
  wire  mem_0_1_R0_data; // @[:anonymous source@346.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@346.4]
  wire [7:0] mem_0_2_W0_addr; // @[:anonymous source@347.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@347.4]
  wire  mem_0_2_W0_data; // @[:anonymous source@347.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@347.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@347.4]
  wire [7:0] mem_0_2_R0_addr; // @[:anonymous source@347.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@347.4]
  wire  mem_0_2_R0_data; // @[:anonymous source@347.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@347.4]
  wire [7:0] mem_0_3_W0_addr; // @[:anonymous source@348.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@348.4]
  wire  mem_0_3_W0_data; // @[:anonymous source@348.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@348.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@348.4]
  wire [7:0] mem_0_3_R0_addr; // @[:anonymous source@348.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@348.4]
  wire  mem_0_3_R0_data; // @[:anonymous source@348.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@348.4]
  wire  R0_data_0_0; // @[:anonymous source@371.4]
  wire  R0_data_0_1; // @[:anonymous source@375.4]
  wire  R0_data_0_2; // @[:anonymous source@379.4]
  wire  R0_data_0_3; // @[:anonymous source@383.4]
  wire [1:0] _GEN_0; // @[:anonymous source@385.4]
  wire [2:0] _GEN_1; // @[:anonymous source@385.4]
  wire [3:0] R0_data_0; // @[:anonymous source@385.4]
  wire [1:0] _GEN_2; // @[:anonymous source@386.4]
  wire [2:0] _GEN_3; // @[:anonymous source@386.4]
  split_hi_us_0_ext mem_0_0 ( // @[:anonymous source@345.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_hi_us_0_ext mem_0_1 ( // @[:anonymous source@346.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_hi_us_0_ext mem_0_2 ( // @[:anonymous source@347.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_hi_us_0_ext mem_0_3 ( // @[:anonymous source@348.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@371.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@375.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@379.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@383.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@385.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@385.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@385.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@386.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@386.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@386.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@350.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@349.4]
  assign mem_0_0_W0_data = W0_data[0]; // @[:anonymous source@351.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@353.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@352.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@370.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@369.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@372.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@355.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@354.4]
  assign mem_0_1_W0_data = W0_data[1]; // @[:anonymous source@356.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@358.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@357.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@374.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@373.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@376.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@360.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@359.4]
  assign mem_0_2_W0_data = W0_data[2]; // @[:anonymous source@361.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@363.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@362.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@378.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@377.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@380.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@365.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@364.4]
  assign mem_0_3_W0_data = W0_data[3]; // @[:anonymous source@366.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@368.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@367.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@382.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@381.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@384.4]
endmodule
module table_0_ext( // @[:anonymous source@388.2]
  input  [7:0]  W0_addr, // @[:anonymous source@389.4]
  input         W0_clk, // @[:anonymous source@390.4]
  input  [47:0] W0_data, // @[:anonymous source@391.4]
  input         W0_en, // @[:anonymous source@392.4]
  input  [3:0]  W0_mask, // @[:anonymous source@393.4]
  input  [7:0]  R0_addr, // @[:anonymous source@394.4]
  input         R0_clk, // @[:anonymous source@395.4]
  output [47:0] R0_data, // @[:anonymous source@396.4]
  input         R0_en // @[:anonymous source@397.4]
);
  wire [7:0] mem_0_0_W0_addr; // @[:anonymous source@399.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@399.4]
  wire [11:0] mem_0_0_W0_data; // @[:anonymous source@399.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@399.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@399.4]
  wire [7:0] mem_0_0_R0_addr; // @[:anonymous source@399.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@399.4]
  wire [11:0] mem_0_0_R0_data; // @[:anonymous source@399.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@399.4]
  wire [7:0] mem_0_1_W0_addr; // @[:anonymous source@400.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@400.4]
  wire [11:0] mem_0_1_W0_data; // @[:anonymous source@400.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@400.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@400.4]
  wire [7:0] mem_0_1_R0_addr; // @[:anonymous source@400.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@400.4]
  wire [11:0] mem_0_1_R0_data; // @[:anonymous source@400.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@400.4]
  wire [7:0] mem_0_2_W0_addr; // @[:anonymous source@401.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@401.4]
  wire [11:0] mem_0_2_W0_data; // @[:anonymous source@401.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@401.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@401.4]
  wire [7:0] mem_0_2_R0_addr; // @[:anonymous source@401.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@401.4]
  wire [11:0] mem_0_2_R0_data; // @[:anonymous source@401.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@401.4]
  wire [7:0] mem_0_3_W0_addr; // @[:anonymous source@402.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@402.4]
  wire [11:0] mem_0_3_W0_data; // @[:anonymous source@402.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@402.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@402.4]
  wire [7:0] mem_0_3_R0_addr; // @[:anonymous source@402.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@402.4]
  wire [11:0] mem_0_3_R0_data; // @[:anonymous source@402.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@402.4]
  wire [11:0] R0_data_0_0; // @[:anonymous source@425.4]
  wire [11:0] R0_data_0_1; // @[:anonymous source@429.4]
  wire [11:0] R0_data_0_2; // @[:anonymous source@433.4]
  wire [11:0] R0_data_0_3; // @[:anonymous source@437.4]
  wire [23:0] _GEN_0; // @[:anonymous source@439.4]
  wire [35:0] _GEN_1; // @[:anonymous source@439.4]
  wire [47:0] R0_data_0; // @[:anonymous source@439.4]
  wire [23:0] _GEN_2; // @[:anonymous source@440.4]
  wire [35:0] _GEN_3; // @[:anonymous source@440.4]
  split_table_0_ext mem_0_0 ( // @[:anonymous source@399.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_table_0_ext mem_0_1 ( // @[:anonymous source@400.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_table_0_ext mem_0_2 ( // @[:anonymous source@401.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_table_0_ext mem_0_3 ( // @[:anonymous source@402.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@425.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@429.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@433.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@437.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@439.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@439.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@439.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@440.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@440.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@440.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@404.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@403.4]
  assign mem_0_0_W0_data = W0_data[11:0]; // @[:anonymous source@405.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@407.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@406.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@424.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@423.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@426.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@409.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@408.4]
  assign mem_0_1_W0_data = W0_data[23:12]; // @[:anonymous source@410.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@412.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@411.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@428.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@427.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@430.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@414.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@413.4]
  assign mem_0_2_W0_data = W0_data[35:24]; // @[:anonymous source@415.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@417.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@416.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@432.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@431.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@434.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@419.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@418.4]
  assign mem_0_3_W0_data = W0_data[47:36]; // @[:anonymous source@420.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@422.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@421.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@436.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@435.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@438.4]
endmodule
module table_1_ext( // @[:anonymous source@442.2]
  input  [6:0]  W0_addr, // @[:anonymous source@443.4]
  input         W0_clk, // @[:anonymous source@444.4]
  input  [51:0] W0_data, // @[:anonymous source@445.4]
  input         W0_en, // @[:anonymous source@446.4]
  input  [3:0]  W0_mask, // @[:anonymous source@447.4]
  input  [6:0]  R0_addr, // @[:anonymous source@448.4]
  input         R0_clk, // @[:anonymous source@449.4]
  output [51:0] R0_data, // @[:anonymous source@450.4]
  input         R0_en // @[:anonymous source@451.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@453.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@453.4]
  wire [12:0] mem_0_0_W0_data; // @[:anonymous source@453.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@453.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@453.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@453.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@453.4]
  wire [12:0] mem_0_0_R0_data; // @[:anonymous source@453.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@453.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@454.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@454.4]
  wire [12:0] mem_0_1_W0_data; // @[:anonymous source@454.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@454.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@454.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@454.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@454.4]
  wire [12:0] mem_0_1_R0_data; // @[:anonymous source@454.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@454.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@455.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@455.4]
  wire [12:0] mem_0_2_W0_data; // @[:anonymous source@455.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@455.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@455.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@455.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@455.4]
  wire [12:0] mem_0_2_R0_data; // @[:anonymous source@455.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@455.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@456.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@456.4]
  wire [12:0] mem_0_3_W0_data; // @[:anonymous source@456.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@456.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@456.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@456.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@456.4]
  wire [12:0] mem_0_3_R0_data; // @[:anonymous source@456.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@456.4]
  wire [12:0] R0_data_0_0; // @[:anonymous source@479.4]
  wire [12:0] R0_data_0_1; // @[:anonymous source@483.4]
  wire [12:0] R0_data_0_2; // @[:anonymous source@487.4]
  wire [12:0] R0_data_0_3; // @[:anonymous source@491.4]
  wire [25:0] _GEN_0; // @[:anonymous source@493.4]
  wire [38:0] _GEN_1; // @[:anonymous source@493.4]
  wire [51:0] R0_data_0; // @[:anonymous source@493.4]
  wire [25:0] _GEN_2; // @[:anonymous source@494.4]
  wire [38:0] _GEN_3; // @[:anonymous source@494.4]
  split_table_1_ext mem_0_0 ( // @[:anonymous source@453.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_table_1_ext mem_0_1 ( // @[:anonymous source@454.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_table_1_ext mem_0_2 ( // @[:anonymous source@455.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_table_1_ext mem_0_3 ( // @[:anonymous source@456.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@479.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@483.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@487.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@491.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@493.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@493.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@493.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@494.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@494.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@494.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@458.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@457.4]
  assign mem_0_0_W0_data = W0_data[12:0]; // @[:anonymous source@459.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@461.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@460.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@478.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@477.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@480.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@463.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@462.4]
  assign mem_0_1_W0_data = W0_data[25:13]; // @[:anonymous source@464.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@466.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@465.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@482.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@481.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@484.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@468.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@467.4]
  assign mem_0_2_W0_data = W0_data[38:26]; // @[:anonymous source@469.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@471.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@470.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@486.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@485.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@488.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@473.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@472.4]
  assign mem_0_3_W0_data = W0_data[51:39]; // @[:anonymous source@474.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@476.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@475.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@490.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@489.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@492.4]
endmodule
module meta_0_ext( // @[:anonymous source@496.2]
  input  [6:0]   W0_addr, // @[:anonymous source@497.4]
  input          W0_clk, // @[:anonymous source@498.4]
  input  [123:0] W0_data, // @[:anonymous source@499.4]
  input          W0_en, // @[:anonymous source@500.4]
  input  [3:0]   W0_mask, // @[:anonymous source@501.4]
  input  [6:0]   R0_addr, // @[:anonymous source@502.4]
  input          R0_clk, // @[:anonymous source@503.4]
  output [123:0] R0_data, // @[:anonymous source@504.4]
  input          R0_en // @[:anonymous source@505.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@507.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@507.4]
  wire [30:0] mem_0_0_W0_data; // @[:anonymous source@507.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@507.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@507.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@507.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@507.4]
  wire [30:0] mem_0_0_R0_data; // @[:anonymous source@507.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@507.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@508.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@508.4]
  wire [30:0] mem_0_1_W0_data; // @[:anonymous source@508.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@508.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@508.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@508.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@508.4]
  wire [30:0] mem_0_1_R0_data; // @[:anonymous source@508.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@508.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@509.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@509.4]
  wire [30:0] mem_0_2_W0_data; // @[:anonymous source@509.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@509.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@509.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@509.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@509.4]
  wire [30:0] mem_0_2_R0_data; // @[:anonymous source@509.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@509.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@510.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@510.4]
  wire [30:0] mem_0_3_W0_data; // @[:anonymous source@510.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@510.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@510.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@510.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@510.4]
  wire [30:0] mem_0_3_R0_data; // @[:anonymous source@510.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@510.4]
  wire [30:0] R0_data_0_0; // @[:anonymous source@533.4]
  wire [30:0] R0_data_0_1; // @[:anonymous source@537.4]
  wire [30:0] R0_data_0_2; // @[:anonymous source@541.4]
  wire [30:0] R0_data_0_3; // @[:anonymous source@545.4]
  wire [61:0] _GEN_0; // @[:anonymous source@547.4]
  wire [92:0] _GEN_1; // @[:anonymous source@547.4]
  wire [123:0] R0_data_0; // @[:anonymous source@547.4]
  wire [61:0] _GEN_2; // @[:anonymous source@548.4]
  wire [92:0] _GEN_3; // @[:anonymous source@548.4]
  split_meta_0_ext mem_0_0 ( // @[:anonymous source@507.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_meta_0_ext mem_0_1 ( // @[:anonymous source@508.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_meta_0_ext mem_0_2 ( // @[:anonymous source@509.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_meta_0_ext mem_0_3 ( // @[:anonymous source@510.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@533.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@537.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@541.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@545.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@547.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@547.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@547.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@548.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@548.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@548.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@512.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@511.4]
  assign mem_0_0_W0_data = W0_data[30:0]; // @[:anonymous source@513.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@515.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@514.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@532.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@531.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@534.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@517.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@516.4]
  assign mem_0_1_W0_data = W0_data[61:31]; // @[:anonymous source@518.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@520.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@519.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@536.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@535.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@538.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@522.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@521.4]
  assign mem_0_2_W0_data = W0_data[92:62]; // @[:anonymous source@523.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@525.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@524.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@540.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@539.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@542.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@527.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@526.4]
  assign mem_0_3_W0_data = W0_data[123:93]; // @[:anonymous source@528.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@530.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@529.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@544.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@543.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@546.4]
endmodule
module btb_0_ext( // @[:anonymous source@550.2]
  input  [6:0]  W0_addr, // @[:anonymous source@551.4]
  input         W0_clk, // @[:anonymous source@552.4]
  input  [55:0] W0_data, // @[:anonymous source@553.4]
  input         W0_en, // @[:anonymous source@554.4]
  input  [3:0]  W0_mask, // @[:anonymous source@555.4]
  input  [6:0]  R0_addr, // @[:anonymous source@556.4]
  input         R0_clk, // @[:anonymous source@557.4]
  output [55:0] R0_data, // @[:anonymous source@558.4]
  input         R0_en // @[:anonymous source@559.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@561.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@561.4]
  wire [13:0] mem_0_0_W0_data; // @[:anonymous source@561.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@561.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@561.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@561.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@561.4]
  wire [13:0] mem_0_0_R0_data; // @[:anonymous source@561.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@561.4]
  wire [6:0] mem_0_1_W0_addr; // @[:anonymous source@562.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@562.4]
  wire [13:0] mem_0_1_W0_data; // @[:anonymous source@562.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@562.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@562.4]
  wire [6:0] mem_0_1_R0_addr; // @[:anonymous source@562.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@562.4]
  wire [13:0] mem_0_1_R0_data; // @[:anonymous source@562.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@562.4]
  wire [6:0] mem_0_2_W0_addr; // @[:anonymous source@563.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@563.4]
  wire [13:0] mem_0_2_W0_data; // @[:anonymous source@563.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@563.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@563.4]
  wire [6:0] mem_0_2_R0_addr; // @[:anonymous source@563.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@563.4]
  wire [13:0] mem_0_2_R0_data; // @[:anonymous source@563.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@563.4]
  wire [6:0] mem_0_3_W0_addr; // @[:anonymous source@564.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@564.4]
  wire [13:0] mem_0_3_W0_data; // @[:anonymous source@564.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@564.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@564.4]
  wire [6:0] mem_0_3_R0_addr; // @[:anonymous source@564.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@564.4]
  wire [13:0] mem_0_3_R0_data; // @[:anonymous source@564.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@564.4]
  wire [13:0] R0_data_0_0; // @[:anonymous source@587.4]
  wire [13:0] R0_data_0_1; // @[:anonymous source@591.4]
  wire [13:0] R0_data_0_2; // @[:anonymous source@595.4]
  wire [13:0] R0_data_0_3; // @[:anonymous source@599.4]
  wire [27:0] _GEN_0; // @[:anonymous source@601.4]
  wire [41:0] _GEN_1; // @[:anonymous source@601.4]
  wire [55:0] R0_data_0; // @[:anonymous source@601.4]
  wire [27:0] _GEN_2; // @[:anonymous source@602.4]
  wire [41:0] _GEN_3; // @[:anonymous source@602.4]
  split_btb_0_ext mem_0_0 ( // @[:anonymous source@561.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_btb_0_ext mem_0_1 ( // @[:anonymous source@562.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_btb_0_ext mem_0_2 ( // @[:anonymous source@563.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_btb_0_ext mem_0_3 ( // @[:anonymous source@564.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@587.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@591.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@595.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@599.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@601.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@601.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@601.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@602.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@602.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@602.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@566.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@565.4]
  assign mem_0_0_W0_data = W0_data[13:0]; // @[:anonymous source@567.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@569.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@568.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@586.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@585.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@588.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@571.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@570.4]
  assign mem_0_1_W0_data = W0_data[27:14]; // @[:anonymous source@572.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@574.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@573.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@590.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@589.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@592.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@576.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@575.4]
  assign mem_0_2_W0_data = W0_data[41:28]; // @[:anonymous source@577.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@579.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@578.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@594.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@593.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@596.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@581.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@580.4]
  assign mem_0_3_W0_data = W0_data[55:42]; // @[:anonymous source@582.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@584.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@583.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@598.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@597.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@600.4]
endmodule
module ebtb_ext( // @[:anonymous source@604.2]
  input  [6:0]  W0_addr, // @[:anonymous source@605.4]
  input         W0_clk, // @[:anonymous source@606.4]
  input  [39:0] W0_data, // @[:anonymous source@607.4]
  input         W0_en, // @[:anonymous source@608.4]
  input  [6:0]  R0_addr, // @[:anonymous source@609.4]
  input         R0_clk, // @[:anonymous source@610.4]
  output [39:0] R0_data, // @[:anonymous source@611.4]
  input         R0_en // @[:anonymous source@612.4]
);
  wire [6:0] mem_0_0_W0_addr; // @[:anonymous source@614.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@614.4]
  wire [39:0] mem_0_0_W0_data; // @[:anonymous source@614.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@614.4]
  wire [6:0] mem_0_0_R0_addr; // @[:anonymous source@614.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@614.4]
  wire [39:0] mem_0_0_R0_data; // @[:anonymous source@614.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@614.4]
  wire [39:0] R0_data_0_0; // @[:anonymous source@621.4]
  wire [39:0] R0_data_0; // @[:anonymous source@623.4]
  split_ebtb_ext mem_0_0 ( // @[:anonymous source@614.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@621.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@623.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@624.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@616.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@615.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@617.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@618.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@620.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@619.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@622.4]
endmodule
module data_ext( // @[:anonymous source@626.2]
  input  [10:0] W0_addr, // @[:anonymous source@627.4]
  input         W0_clk, // @[:anonymous source@628.4]
  input  [7:0]  W0_data, // @[:anonymous source@629.4]
  input         W0_en, // @[:anonymous source@630.4]
  input  [3:0]  W0_mask, // @[:anonymous source@631.4]
  input  [10:0] R0_addr, // @[:anonymous source@632.4]
  input         R0_clk, // @[:anonymous source@633.4]
  output [7:0]  R0_data, // @[:anonymous source@634.4]
  input         R0_en // @[:anonymous source@635.4]
);
  wire [10:0] mem_0_0_W0_addr; // @[:anonymous source@637.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@637.4]
  wire [1:0] mem_0_0_W0_data; // @[:anonymous source@637.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@637.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@637.4]
  wire [10:0] mem_0_0_R0_addr; // @[:anonymous source@637.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@637.4]
  wire [1:0] mem_0_0_R0_data; // @[:anonymous source@637.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@637.4]
  wire [10:0] mem_0_1_W0_addr; // @[:anonymous source@638.4]
  wire  mem_0_1_W0_clk; // @[:anonymous source@638.4]
  wire [1:0] mem_0_1_W0_data; // @[:anonymous source@638.4]
  wire  mem_0_1_W0_en; // @[:anonymous source@638.4]
  wire  mem_0_1_W0_mask; // @[:anonymous source@638.4]
  wire [10:0] mem_0_1_R0_addr; // @[:anonymous source@638.4]
  wire  mem_0_1_R0_clk; // @[:anonymous source@638.4]
  wire [1:0] mem_0_1_R0_data; // @[:anonymous source@638.4]
  wire  mem_0_1_R0_en; // @[:anonymous source@638.4]
  wire [10:0] mem_0_2_W0_addr; // @[:anonymous source@639.4]
  wire  mem_0_2_W0_clk; // @[:anonymous source@639.4]
  wire [1:0] mem_0_2_W0_data; // @[:anonymous source@639.4]
  wire  mem_0_2_W0_en; // @[:anonymous source@639.4]
  wire  mem_0_2_W0_mask; // @[:anonymous source@639.4]
  wire [10:0] mem_0_2_R0_addr; // @[:anonymous source@639.4]
  wire  mem_0_2_R0_clk; // @[:anonymous source@639.4]
  wire [1:0] mem_0_2_R0_data; // @[:anonymous source@639.4]
  wire  mem_0_2_R0_en; // @[:anonymous source@639.4]
  wire [10:0] mem_0_3_W0_addr; // @[:anonymous source@640.4]
  wire  mem_0_3_W0_clk; // @[:anonymous source@640.4]
  wire [1:0] mem_0_3_W0_data; // @[:anonymous source@640.4]
  wire  mem_0_3_W0_en; // @[:anonymous source@640.4]
  wire  mem_0_3_W0_mask; // @[:anonymous source@640.4]
  wire [10:0] mem_0_3_R0_addr; // @[:anonymous source@640.4]
  wire  mem_0_3_R0_clk; // @[:anonymous source@640.4]
  wire [1:0] mem_0_3_R0_data; // @[:anonymous source@640.4]
  wire  mem_0_3_R0_en; // @[:anonymous source@640.4]
  wire [1:0] R0_data_0_0; // @[:anonymous source@663.4]
  wire [1:0] R0_data_0_1; // @[:anonymous source@667.4]
  wire [1:0] R0_data_0_2; // @[:anonymous source@671.4]
  wire [1:0] R0_data_0_3; // @[:anonymous source@675.4]
  wire [3:0] _GEN_0; // @[:anonymous source@677.4]
  wire [5:0] _GEN_1; // @[:anonymous source@677.4]
  wire [7:0] R0_data_0; // @[:anonymous source@677.4]
  wire [3:0] _GEN_2; // @[:anonymous source@678.4]
  wire [5:0] _GEN_3; // @[:anonymous source@678.4]
  split_data_ext mem_0_0 ( // @[:anonymous source@637.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  split_data_ext mem_0_1 ( // @[:anonymous source@638.4]
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask),
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en)
  );
  split_data_ext mem_0_2 ( // @[:anonymous source@639.4]
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask),
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en)
  );
  split_data_ext mem_0_3 ( // @[:anonymous source@640.4]
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask),
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@663.4]
  assign R0_data_0_1 = mem_0_1_R0_data; // @[:anonymous source@667.4]
  assign R0_data_0_2 = mem_0_2_R0_data; // @[:anonymous source@671.4]
  assign R0_data_0_3 = mem_0_3_R0_data; // @[:anonymous source@675.4]
  assign _GEN_0 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@677.4]
  assign _GEN_1 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@677.4]
  assign R0_data_0 = {R0_data_0_3,R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@677.4]
  assign _GEN_2 = {R0_data_0_1,R0_data_0_0}; // @[:anonymous source@678.4]
  assign _GEN_3 = {R0_data_0_2,R0_data_0_1,R0_data_0_0}; // @[:anonymous source@678.4]
  assign R0_data = {R0_data_0_3,_GEN_1}; // @[:anonymous source@678.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@642.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@641.4]
  assign mem_0_0_W0_data = W0_data[1:0]; // @[:anonymous source@643.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@645.4]
  assign mem_0_0_W0_mask = W0_mask[0]; // @[:anonymous source@644.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@662.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@661.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@664.4]
  assign mem_0_1_W0_addr = W0_addr; // @[:anonymous source@647.4]
  assign mem_0_1_W0_clk = W0_clk; // @[:anonymous source@646.4]
  assign mem_0_1_W0_data = W0_data[3:2]; // @[:anonymous source@648.4]
  assign mem_0_1_W0_en = W0_en; // @[:anonymous source@650.4]
  assign mem_0_1_W0_mask = W0_mask[1]; // @[:anonymous source@649.4]
  assign mem_0_1_R0_addr = R0_addr; // @[:anonymous source@666.4]
  assign mem_0_1_R0_clk = R0_clk; // @[:anonymous source@665.4]
  assign mem_0_1_R0_en = R0_en; // @[:anonymous source@668.4]
  assign mem_0_2_W0_addr = W0_addr; // @[:anonymous source@652.4]
  assign mem_0_2_W0_clk = W0_clk; // @[:anonymous source@651.4]
  assign mem_0_2_W0_data = W0_data[5:4]; // @[:anonymous source@653.4]
  assign mem_0_2_W0_en = W0_en; // @[:anonymous source@655.4]
  assign mem_0_2_W0_mask = W0_mask[2]; // @[:anonymous source@654.4]
  assign mem_0_2_R0_addr = R0_addr; // @[:anonymous source@670.4]
  assign mem_0_2_R0_clk = R0_clk; // @[:anonymous source@669.4]
  assign mem_0_2_R0_en = R0_en; // @[:anonymous source@672.4]
  assign mem_0_3_W0_addr = W0_addr; // @[:anonymous source@657.4]
  assign mem_0_3_W0_clk = W0_clk; // @[:anonymous source@656.4]
  assign mem_0_3_W0_data = W0_data[7:6]; // @[:anonymous source@658.4]
  assign mem_0_3_W0_en = W0_en; // @[:anonymous source@660.4]
  assign mem_0_3_W0_mask = W0_mask[3]; // @[:anonymous source@659.4]
  assign mem_0_3_R0_addr = R0_addr; // @[:anonymous source@674.4]
  assign mem_0_3_R0_clk = R0_clk; // @[:anonymous source@673.4]
  assign mem_0_3_R0_en = R0_en; // @[:anonymous source@676.4]
endmodule
module meta_ext( // @[:anonymous source@680.2]
  input  [3:0]   W0_addr, // @[:anonymous source@681.4]
  input          W0_clk, // @[:anonymous source@682.4]
  input  [119:0] W0_data, // @[:anonymous source@683.4]
  input          W0_en, // @[:anonymous source@684.4]
  input  [3:0]   R0_addr, // @[:anonymous source@685.4]
  input          R0_clk, // @[:anonymous source@686.4]
  output [119:0] R0_data, // @[:anonymous source@687.4]
  input          R0_en // @[:anonymous source@688.4]
);
  wire [3:0] mem_0_0_W0_addr; // @[:anonymous source@690.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@690.4]
  wire [119:0] mem_0_0_W0_data; // @[:anonymous source@690.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@690.4]
  wire [3:0] mem_0_0_R0_addr; // @[:anonymous source@690.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@690.4]
  wire [119:0] mem_0_0_R0_data; // @[:anonymous source@690.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@690.4]
  wire [119:0] R0_data_0_0; // @[:anonymous source@697.4]
  wire [119:0] R0_data_0; // @[:anonymous source@699.4]
  split_meta_ext mem_0_0 ( // @[:anonymous source@690.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@697.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@699.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@700.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@692.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@691.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@693.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@694.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@696.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@695.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@698.4]
endmodule
module ghist_0_ext( // @[:anonymous source@702.2]
  input  [3:0]  W0_addr, // @[:anonymous source@703.4]
  input         W0_clk, // @[:anonymous source@704.4]
  input  [71:0] W0_data, // @[:anonymous source@705.4]
  input         W0_en, // @[:anonymous source@706.4]
  input  [3:0]  R0_addr, // @[:anonymous source@707.4]
  input         R0_clk, // @[:anonymous source@708.4]
  output [71:0] R0_data, // @[:anonymous source@709.4]
  input         R0_en // @[:anonymous source@710.4]
);
  wire [3:0] mem_0_0_W0_addr; // @[:anonymous source@712.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@712.4]
  wire [71:0] mem_0_0_W0_data; // @[:anonymous source@712.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@712.4]
  wire [3:0] mem_0_0_R0_addr; // @[:anonymous source@712.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@712.4]
  wire [71:0] mem_0_0_R0_data; // @[:anonymous source@712.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@712.4]
  wire [71:0] R0_data_0_0; // @[:anonymous source@719.4]
  wire [71:0] R0_data_0; // @[:anonymous source@721.4]
  split_ghist_0_ext mem_0_0 ( // @[:anonymous source@712.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@719.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@721.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@722.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@714.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@713.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@715.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@716.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@718.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@717.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@720.4]
endmodule
module rob_debug_inst_mem_ext( // @[:anonymous source@724.2]
  input  [4:0]  W0_addr, // @[:anonymous source@725.4]
  input         W0_clk, // @[:anonymous source@726.4]
  input  [31:0] W0_data, // @[:anonymous source@727.4]
  input         W0_en, // @[:anonymous source@728.4]
  input         W0_mask, // @[:anonymous source@729.4]
  input  [4:0]  R0_addr, // @[:anonymous source@730.4]
  input         R0_clk, // @[:anonymous source@731.4]
  output [31:0] R0_data, // @[:anonymous source@732.4]
  input         R0_en // @[:anonymous source@733.4]
);
  wire [4:0] mem_0_0_W0_addr; // @[:anonymous source@735.4]
  wire  mem_0_0_W0_clk; // @[:anonymous source@735.4]
  wire [31:0] mem_0_0_W0_data; // @[:anonymous source@735.4]
  wire  mem_0_0_W0_en; // @[:anonymous source@735.4]
  wire  mem_0_0_W0_mask; // @[:anonymous source@735.4]
  wire [4:0] mem_0_0_R0_addr; // @[:anonymous source@735.4]
  wire  mem_0_0_R0_clk; // @[:anonymous source@735.4]
  wire [31:0] mem_0_0_R0_data; // @[:anonymous source@735.4]
  wire  mem_0_0_R0_en; // @[:anonymous source@735.4]
  wire [31:0] R0_data_0_0; // @[:anonymous source@743.4]
  wire [31:0] R0_data_0; // @[:anonymous source@745.4]
  split_rob_debug_inst_mem_ext mem_0_0 ( // @[:anonymous source@735.4]
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask),
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en)
  );
  assign R0_data_0_0 = mem_0_0_R0_data; // @[:anonymous source@743.4]
  assign R0_data_0 = R0_data_0_0; // @[:anonymous source@745.4]
  assign R0_data = mem_0_0_R0_data; // @[:anonymous source@746.4]
  assign mem_0_0_W0_addr = W0_addr; // @[:anonymous source@737.4]
  assign mem_0_0_W0_clk = W0_clk; // @[:anonymous source@736.4]
  assign mem_0_0_W0_data = W0_data; // @[:anonymous source@738.4]
  assign mem_0_0_W0_en = W0_en; // @[:anonymous source@740.4]
  assign mem_0_0_W0_mask = W0_mask; // @[:anonymous source@739.4]
  assign mem_0_0_R0_addr = R0_addr; // @[:anonymous source@742.4]
  assign mem_0_0_R0_clk = R0_clk; // @[:anonymous source@741.4]
  assign mem_0_0_R0_en = R0_en; // @[:anonymous source@744.4]
endmodule
module l2_tlb_ram_ext( // @[:anonymous source@748.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@749.4]
  input         RW0_clk, // @[:anonymous source@750.4]
  input  [43:0] RW0_wdata, // @[:anonymous source@751.4]
  output [43:0] RW0_rdata, // @[:anonymous source@752.4]
  input         RW0_en, // @[:anonymous source@753.4]
  input         RW0_wmode // @[:anonymous source@754.4]
);
  wire [9:0] mem_0_0_RW0_addr; // @[:anonymous source@756.4]
  wire  mem_0_0_RW0_clk; // @[:anonymous source@756.4]
  wire [43:0] mem_0_0_RW0_wdata; // @[:anonymous source@756.4]
  wire [43:0] mem_0_0_RW0_rdata; // @[:anonymous source@756.4]
  wire  mem_0_0_RW0_en; // @[:anonymous source@756.4]
  wire  mem_0_0_RW0_wmode; // @[:anonymous source@756.4]
  wire [43:0] RW0_rdata_0_0; // @[:anonymous source@759.4]
  wire [43:0] RW0_rdata_0; // @[:anonymous source@763.4]
  split_l2_tlb_ram_ext mem_0_0 ( // @[:anonymous source@756.4]
    .RW0_addr(mem_0_0_RW0_addr),
    .RW0_clk(mem_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_RW0_rdata),
    .RW0_en(mem_0_0_RW0_en),
    .RW0_wmode(mem_0_0_RW0_wmode)
  );
  assign RW0_rdata_0_0 = mem_0_0_RW0_rdata; // @[:anonymous source@759.4]
  assign RW0_rdata_0 = RW0_rdata_0_0; // @[:anonymous source@763.4]
  assign RW0_rdata = mem_0_0_RW0_rdata; // @[:anonymous source@764.4]
  assign mem_0_0_RW0_addr = RW0_addr; // @[:anonymous source@758.4]
  assign mem_0_0_RW0_clk = RW0_clk; // @[:anonymous source@757.4]
  assign mem_0_0_RW0_wdata = RW0_wdata; // @[:anonymous source@760.4]
  assign mem_0_0_RW0_en = RW0_en; // @[:anonymous source@762.4]
  assign mem_0_0_RW0_wmode = RW0_wmode; // @[:anonymous source@761.4]
endmodule
module split_cc_dir_ext( // @[:anonymous source@766.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@767.4]
  input         RW0_clk, // @[:anonymous source@768.4]
  input  [15:0] RW0_wdata, // @[:anonymous source@769.4]
  output [15:0] RW0_rdata, // @[:anonymous source@770.4]
  input         RW0_en, // @[:anonymous source@771.4]
  input         RW0_wmode, // @[:anonymous source@772.4]
  input         RW0_wmask // @[:anonymous source@773.4]
);
  reg [15:0] ram [0:1023]; // @[:anonymous source@775.4]
  reg [31:0] _RAND_0;
  wire [15:0] ram_RW_0_r_data; // @[:anonymous source@775.4]
  wire [9:0] ram_RW_0_r_addr; // @[:anonymous source@775.4]
  wire [15:0] ram_RW_0_w_data; // @[:anonymous source@775.4]
  wire [9:0] ram_RW_0_w_addr; // @[:anonymous source@775.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@775.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@775.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [9:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@775.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@787.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[15:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@775.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_cc_banks_0_ext( // @[:anonymous source@790.2]
  input  [13:0] RW0_addr, // @[:anonymous source@791.4]
  input         RW0_clk, // @[:anonymous source@792.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@793.4]
  output [63:0] RW0_rdata, // @[:anonymous source@794.4]
  input         RW0_en, // @[:anonymous source@795.4]
  input         RW0_wmode // @[:anonymous source@796.4]
);
  reg [63:0] ram [0:16383]; // @[:anonymous source@798.4]
  reg [63:0] _RAND_0;
  wire [63:0] ram_RW_0_r_data; // @[:anonymous source@798.4]
  wire [13:0] ram_RW_0_r_addr; // @[:anonymous source@798.4]
  wire [63:0] ram_RW_0_w_data; // @[:anonymous source@798.4]
  wire [13:0] ram_RW_0_w_addr; // @[:anonymous source@798.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@798.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@798.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [13:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@798.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@810.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16384; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@798.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_tag_array_ext( // @[:anonymous source@813.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@814.4]
  input         RW0_clk, // @[:anonymous source@815.4]
  input  [21:0] RW0_wdata, // @[:anonymous source@816.4]
  output [21:0] RW0_rdata, // @[:anonymous source@817.4]
  input         RW0_en, // @[:anonymous source@818.4]
  input         RW0_wmode, // @[:anonymous source@819.4]
  input         RW0_wmask // @[:anonymous source@820.4]
);
  reg [21:0] ram [0:63]; // @[:anonymous source@822.4]
  reg [31:0] _RAND_0;
  wire [21:0] ram_RW_0_r_data; // @[:anonymous source@822.4]
  wire [5:0] ram_RW_0_r_addr; // @[:anonymous source@822.4]
  wire [21:0] ram_RW_0_w_data; // @[:anonymous source@822.4]
  wire [5:0] ram_RW_0_w_addr; // @[:anonymous source@822.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@822.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@822.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@822.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@834.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[21:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@822.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_array_0_0_ext( // @[:anonymous source@837.2]
  input  [8:0]  W0_addr, // @[:anonymous source@838.4]
  input         W0_clk, // @[:anonymous source@839.4]
  input  [63:0] W0_data, // @[:anonymous source@840.4]
  input         W0_en, // @[:anonymous source@841.4]
  input         W0_mask, // @[:anonymous source@842.4]
  input  [8:0]  R0_addr, // @[:anonymous source@843.4]
  input         R0_clk, // @[:anonymous source@844.4]
  output [63:0] R0_data, // @[:anonymous source@845.4]
  input         R0_en // @[:anonymous source@846.4]
);
  reg [63:0] ram [0:511]; // @[:anonymous source@848.4]
  reg [63:0] _RAND_0;
  wire [63:0] ram_R_0_data; // @[:anonymous source@848.4]
  wire [8:0] ram_R_0_addr; // @[:anonymous source@848.4]
  wire [63:0] ram_W_0_data; // @[:anonymous source@848.4]
  wire [8:0] ram_W_0_addr; // @[:anonymous source@848.4]
  wire  ram_W_0_mask; // @[:anonymous source@848.4]
  wire  ram_W_0_en; // @[:anonymous source@848.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [8:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@848.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@859.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@848.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_tag_array_0_ext( // @[:anonymous source@866.2]
  input  [5:0]  RW0_addr, // @[:anonymous source@867.4]
  input         RW0_clk, // @[:anonymous source@868.4]
  input  [19:0] RW0_wdata, // @[:anonymous source@869.4]
  output [19:0] RW0_rdata, // @[:anonymous source@870.4]
  input         RW0_en, // @[:anonymous source@871.4]
  input         RW0_wmode, // @[:anonymous source@872.4]
  input         RW0_wmask // @[:anonymous source@873.4]
);
  reg [19:0] ram [0:63]; // @[:anonymous source@875.4]
  reg [31:0] _RAND_0;
  wire [19:0] ram_RW_0_r_data; // @[:anonymous source@875.4]
  wire [5:0] ram_RW_0_r_addr; // @[:anonymous source@875.4]
  wire [19:0] ram_RW_0_w_data; // @[:anonymous source@875.4]
  wire [5:0] ram_RW_0_w_addr; // @[:anonymous source@875.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@875.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@875.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [5:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@875.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@887.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    ram[initvar] = _RAND_0[19:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[5:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@875.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_dataArrayWay_0_ext( // @[:anonymous source@890.2]
  input  [8:0]  RW0_addr, // @[:anonymous source@891.4]
  input         RW0_clk, // @[:anonymous source@892.4]
  input  [63:0] RW0_wdata, // @[:anonymous source@893.4]
  output [63:0] RW0_rdata, // @[:anonymous source@894.4]
  input         RW0_en, // @[:anonymous source@895.4]
  input         RW0_wmode // @[:anonymous source@896.4]
);
  reg [63:0] ram [0:511]; // @[:anonymous source@898.4]
  reg [63:0] _RAND_0;
  wire [63:0] ram_RW_0_r_data; // @[:anonymous source@898.4]
  wire [8:0] ram_RW_0_r_addr; // @[:anonymous source@898.4]
  wire [63:0] ram_RW_0_w_data; // @[:anonymous source@898.4]
  wire [8:0] ram_RW_0_w_addr; // @[:anonymous source@898.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@898.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@898.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [8:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@898.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@910.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    ram[initvar] = _RAND_0[63:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[8:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@898.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
module split_hi_us_ext( // @[:anonymous source@913.2]
  input  [6:0] W0_addr, // @[:anonymous source@914.4]
  input        W0_clk, // @[:anonymous source@915.4]
  input        W0_data, // @[:anonymous source@916.4]
  input        W0_en, // @[:anonymous source@917.4]
  input        W0_mask, // @[:anonymous source@918.4]
  input  [6:0] R0_addr, // @[:anonymous source@919.4]
  input        R0_clk, // @[:anonymous source@920.4]
  output       R0_data, // @[:anonymous source@921.4]
  input        R0_en // @[:anonymous source@922.4]
);
  reg  ram [0:127]; // @[:anonymous source@924.4]
  reg [31:0] _RAND_0;
  wire  ram_R_0_data; // @[:anonymous source@924.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@924.4]
  wire  ram_W_0_data; // @[:anonymous source@924.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@924.4]
  wire  ram_W_0_mask; // @[:anonymous source@924.4]
  wire  ram_W_0_en; // @[:anonymous source@924.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@924.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@935.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@924.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_table_ext( // @[:anonymous source@942.2]
  input  [6:0]  W0_addr, // @[:anonymous source@943.4]
  input         W0_clk, // @[:anonymous source@944.4]
  input  [10:0] W0_data, // @[:anonymous source@945.4]
  input         W0_en, // @[:anonymous source@946.4]
  input         W0_mask, // @[:anonymous source@947.4]
  input  [6:0]  R0_addr, // @[:anonymous source@948.4]
  input         R0_clk, // @[:anonymous source@949.4]
  output [10:0] R0_data, // @[:anonymous source@950.4]
  input         R0_en // @[:anonymous source@951.4]
);
  reg [10:0] ram [0:127]; // @[:anonymous source@953.4]
  reg [31:0] _RAND_0;
  wire [10:0] ram_R_0_data; // @[:anonymous source@953.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@953.4]
  wire [10:0] ram_W_0_data; // @[:anonymous source@953.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@953.4]
  wire  ram_W_0_mask; // @[:anonymous source@953.4]
  wire  ram_W_0_en; // @[:anonymous source@953.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@953.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@964.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[10:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@953.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_hi_us_0_ext( // @[:anonymous source@971.2]
  input  [7:0] W0_addr, // @[:anonymous source@972.4]
  input        W0_clk, // @[:anonymous source@973.4]
  input        W0_data, // @[:anonymous source@974.4]
  input        W0_en, // @[:anonymous source@975.4]
  input        W0_mask, // @[:anonymous source@976.4]
  input  [7:0] R0_addr, // @[:anonymous source@977.4]
  input        R0_clk, // @[:anonymous source@978.4]
  output       R0_data, // @[:anonymous source@979.4]
  input        R0_en // @[:anonymous source@980.4]
);
  reg  ram [0:255]; // @[:anonymous source@982.4]
  reg [31:0] _RAND_0;
  wire  ram_R_0_data; // @[:anonymous source@982.4]
  wire [7:0] ram_R_0_addr; // @[:anonymous source@982.4]
  wire  ram_W_0_data; // @[:anonymous source@982.4]
  wire [7:0] ram_W_0_addr; // @[:anonymous source@982.4]
  wire  ram_W_0_mask; // @[:anonymous source@982.4]
  wire  ram_W_0_en; // @[:anonymous source@982.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@982.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@993.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@982.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_table_0_ext( // @[:anonymous source@1000.2]
  input  [7:0]  W0_addr, // @[:anonymous source@1001.4]
  input         W0_clk, // @[:anonymous source@1002.4]
  input  [11:0] W0_data, // @[:anonymous source@1003.4]
  input         W0_en, // @[:anonymous source@1004.4]
  input         W0_mask, // @[:anonymous source@1005.4]
  input  [7:0]  R0_addr, // @[:anonymous source@1006.4]
  input         R0_clk, // @[:anonymous source@1007.4]
  output [11:0] R0_data, // @[:anonymous source@1008.4]
  input         R0_en // @[:anonymous source@1009.4]
);
  reg [11:0] ram [0:255]; // @[:anonymous source@1011.4]
  reg [31:0] _RAND_0;
  wire [11:0] ram_R_0_data; // @[:anonymous source@1011.4]
  wire [7:0] ram_R_0_addr; // @[:anonymous source@1011.4]
  wire [11:0] ram_W_0_data; // @[:anonymous source@1011.4]
  wire [7:0] ram_W_0_addr; // @[:anonymous source@1011.4]
  wire  ram_W_0_mask; // @[:anonymous source@1011.4]
  wire  ram_W_0_en; // @[:anonymous source@1011.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [7:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1011.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1022.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    ram[initvar] = _RAND_0[11:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1011.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_table_1_ext( // @[:anonymous source@1029.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1030.4]
  input         W0_clk, // @[:anonymous source@1031.4]
  input  [12:0] W0_data, // @[:anonymous source@1032.4]
  input         W0_en, // @[:anonymous source@1033.4]
  input         W0_mask, // @[:anonymous source@1034.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1035.4]
  input         R0_clk, // @[:anonymous source@1036.4]
  output [12:0] R0_data, // @[:anonymous source@1037.4]
  input         R0_en // @[:anonymous source@1038.4]
);
  reg [12:0] ram [0:127]; // @[:anonymous source@1040.4]
  reg [31:0] _RAND_0;
  wire [12:0] ram_R_0_data; // @[:anonymous source@1040.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1040.4]
  wire [12:0] ram_W_0_data; // @[:anonymous source@1040.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1040.4]
  wire  ram_W_0_mask; // @[:anonymous source@1040.4]
  wire  ram_W_0_en; // @[:anonymous source@1040.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1040.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1051.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[12:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1040.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_meta_0_ext( // @[:anonymous source@1058.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1059.4]
  input         W0_clk, // @[:anonymous source@1060.4]
  input  [30:0] W0_data, // @[:anonymous source@1061.4]
  input         W0_en, // @[:anonymous source@1062.4]
  input         W0_mask, // @[:anonymous source@1063.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1064.4]
  input         R0_clk, // @[:anonymous source@1065.4]
  output [30:0] R0_data, // @[:anonymous source@1066.4]
  input         R0_en // @[:anonymous source@1067.4]
);
  reg [30:0] ram [0:127]; // @[:anonymous source@1069.4]
  reg [31:0] _RAND_0;
  wire [30:0] ram_R_0_data; // @[:anonymous source@1069.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1069.4]
  wire [30:0] ram_W_0_data; // @[:anonymous source@1069.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1069.4]
  wire  ram_W_0_mask; // @[:anonymous source@1069.4]
  wire  ram_W_0_en; // @[:anonymous source@1069.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1069.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1080.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[30:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1069.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_btb_0_ext( // @[:anonymous source@1087.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1088.4]
  input         W0_clk, // @[:anonymous source@1089.4]
  input  [13:0] W0_data, // @[:anonymous source@1090.4]
  input         W0_en, // @[:anonymous source@1091.4]
  input         W0_mask, // @[:anonymous source@1092.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1093.4]
  input         R0_clk, // @[:anonymous source@1094.4]
  output [13:0] R0_data, // @[:anonymous source@1095.4]
  input         R0_en // @[:anonymous source@1096.4]
);
  reg [13:0] ram [0:127]; // @[:anonymous source@1098.4]
  reg [31:0] _RAND_0;
  wire [13:0] ram_R_0_data; // @[:anonymous source@1098.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1098.4]
  wire [13:0] ram_W_0_data; // @[:anonymous source@1098.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1098.4]
  wire  ram_W_0_mask; // @[:anonymous source@1098.4]
  wire  ram_W_0_en; // @[:anonymous source@1098.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1098.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1109.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[13:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1098.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_ebtb_ext( // @[:anonymous source@1116.2]
  input  [6:0]  W0_addr, // @[:anonymous source@1117.4]
  input         W0_clk, // @[:anonymous source@1118.4]
  input  [39:0] W0_data, // @[:anonymous source@1119.4]
  input         W0_en, // @[:anonymous source@1120.4]
  input  [6:0]  R0_addr, // @[:anonymous source@1121.4]
  input         R0_clk, // @[:anonymous source@1122.4]
  output [39:0] R0_data, // @[:anonymous source@1123.4]
  input         R0_en // @[:anonymous source@1124.4]
);
  reg [39:0] ram [0:127]; // @[:anonymous source@1126.4]
  reg [63:0] _RAND_0;
  wire [39:0] ram_R_0_data; // @[:anonymous source@1126.4]
  wire [6:0] ram_R_0_addr; // @[:anonymous source@1126.4]
  wire [39:0] ram_W_0_data; // @[:anonymous source@1126.4]
  wire [6:0] ram_W_0_addr; // @[:anonymous source@1126.4]
  wire  ram_W_0_mask; // @[:anonymous source@1126.4]
  wire  ram_W_0_en; // @[:anonymous source@1126.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [6:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1126.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = 1'h1;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1137.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    ram[initvar] = _RAND_0[39:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1126.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_data_ext( // @[:anonymous source@1144.2]
  input  [10:0] W0_addr, // @[:anonymous source@1145.4]
  input         W0_clk, // @[:anonymous source@1146.4]
  input  [1:0]  W0_data, // @[:anonymous source@1147.4]
  input         W0_en, // @[:anonymous source@1148.4]
  input         W0_mask, // @[:anonymous source@1149.4]
  input  [10:0] R0_addr, // @[:anonymous source@1150.4]
  input         R0_clk, // @[:anonymous source@1151.4]
  output [1:0]  R0_data, // @[:anonymous source@1152.4]
  input         R0_en // @[:anonymous source@1153.4]
);
  reg [1:0] ram [0:2047]; // @[:anonymous source@1155.4]
  reg [31:0] _RAND_0;
  wire [1:0] ram_R_0_data; // @[:anonymous source@1155.4]
  wire [10:0] ram_R_0_addr; // @[:anonymous source@1155.4]
  wire [1:0] ram_W_0_data; // @[:anonymous source@1155.4]
  wire [10:0] ram_W_0_addr; // @[:anonymous source@1155.4]
  wire  ram_W_0_mask; // @[:anonymous source@1155.4]
  wire  ram_W_0_en; // @[:anonymous source@1155.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [10:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1155.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1166.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    ram[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[10:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1155.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_meta_ext( // @[:anonymous source@1173.2]
  input  [3:0]   W0_addr, // @[:anonymous source@1174.4]
  input          W0_clk, // @[:anonymous source@1175.4]
  input  [119:0] W0_data, // @[:anonymous source@1176.4]
  input          W0_en, // @[:anonymous source@1177.4]
  input  [3:0]   R0_addr, // @[:anonymous source@1178.4]
  input          R0_clk, // @[:anonymous source@1179.4]
  output [119:0] R0_data, // @[:anonymous source@1180.4]
  input          R0_en // @[:anonymous source@1181.4]
);
  reg [119:0] ram [0:15]; // @[:anonymous source@1183.4]
  reg [127:0] _RAND_0;
  wire [119:0] ram_R_0_data; // @[:anonymous source@1183.4]
  wire [3:0] ram_R_0_addr; // @[:anonymous source@1183.4]
  wire [119:0] ram_W_0_data; // @[:anonymous source@1183.4]
  wire [3:0] ram_W_0_addr; // @[:anonymous source@1183.4]
  wire  ram_W_0_mask; // @[:anonymous source@1183.4]
  wire  ram_W_0_en; // @[:anonymous source@1183.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [3:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1183.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = 1'h1;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1194.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {4{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[119:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1183.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_ghist_0_ext( // @[:anonymous source@1201.2]
  input  [3:0]  W0_addr, // @[:anonymous source@1202.4]
  input         W0_clk, // @[:anonymous source@1203.4]
  input  [71:0] W0_data, // @[:anonymous source@1204.4]
  input         W0_en, // @[:anonymous source@1205.4]
  input  [3:0]  R0_addr, // @[:anonymous source@1206.4]
  input         R0_clk, // @[:anonymous source@1207.4]
  output [71:0] R0_data, // @[:anonymous source@1208.4]
  input         R0_en // @[:anonymous source@1209.4]
);
  reg [71:0] ram [0:15]; // @[:anonymous source@1211.4]
  reg [95:0] _RAND_0;
  wire [71:0] ram_R_0_data; // @[:anonymous source@1211.4]
  wire [3:0] ram_R_0_addr; // @[:anonymous source@1211.4]
  wire [71:0] ram_W_0_data; // @[:anonymous source@1211.4]
  wire [3:0] ram_W_0_addr; // @[:anonymous source@1211.4]
  wire  ram_W_0_mask; // @[:anonymous source@1211.4]
  wire  ram_W_0_en; // @[:anonymous source@1211.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [3:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1211.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = 1'h1;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1222.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {3{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ram[initvar] = _RAND_0[71:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1211.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_rob_debug_inst_mem_ext( // @[:anonymous source@1229.2]
  input  [4:0]  W0_addr, // @[:anonymous source@1230.4]
  input         W0_clk, // @[:anonymous source@1231.4]
  input  [31:0] W0_data, // @[:anonymous source@1232.4]
  input         W0_en, // @[:anonymous source@1233.4]
  input         W0_mask, // @[:anonymous source@1234.4]
  input  [4:0]  R0_addr, // @[:anonymous source@1235.4]
  input         R0_clk, // @[:anonymous source@1236.4]
  output [31:0] R0_data, // @[:anonymous source@1237.4]
  input         R0_en // @[:anonymous source@1238.4]
);
  reg [31:0] ram [0:31]; // @[:anonymous source@1240.4]
  reg [31:0] _RAND_0;
  wire [31:0] ram_R_0_data; // @[:anonymous source@1240.4]
  wire [4:0] ram_R_0_addr; // @[:anonymous source@1240.4]
  wire [31:0] ram_W_0_data; // @[:anonymous source@1240.4]
  wire [4:0] ram_W_0_addr; // @[:anonymous source@1240.4]
  wire  ram_W_0_mask; // @[:anonymous source@1240.4]
  wire  ram_W_0_en; // @[:anonymous source@1240.4]
  reg  ram_R_0_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [4:0] ram_R_0_addr_pipe_0;
  reg [31:0] _RAND_2;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr]; // @[:anonymous source@1240.4]
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data; // @[:anonymous source@1251.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge W0_clk) begin
    if(ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data; // @[:anonymous source@1240.4]
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
endmodule
module split_l2_tlb_ram_ext( // @[:anonymous source@1258.2]
  input  [9:0]  RW0_addr, // @[:anonymous source@1259.4]
  input         RW0_clk, // @[:anonymous source@1260.4]
  input  [43:0] RW0_wdata, // @[:anonymous source@1261.4]
  output [43:0] RW0_rdata, // @[:anonymous source@1262.4]
  input         RW0_en, // @[:anonymous source@1263.4]
  input         RW0_wmode // @[:anonymous source@1264.4]
);
  reg [43:0] ram [0:1023]; // @[:anonymous source@1266.4]
  reg [63:0] _RAND_0;
  wire [43:0] ram_RW_0_r_data; // @[:anonymous source@1266.4]
  wire [9:0] ram_RW_0_r_addr; // @[:anonymous source@1266.4]
  wire [43:0] ram_RW_0_w_data; // @[:anonymous source@1266.4]
  wire [9:0] ram_RW_0_w_addr; // @[:anonymous source@1266.4]
  wire  ram_RW_0_w_mask; // @[:anonymous source@1266.4]
  wire  ram_RW_0_w_en; // @[:anonymous source@1266.4]
  reg  ram_RW_0_r_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [9:0] ram_RW_0_r_addr_pipe_0;
  reg [31:0] _RAND_2;
  wire  _GEN_0;
  wire  _GEN_1;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr]; // @[:anonymous source@1266.4]
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = 1'h1;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data; // @[:anonymous source@1278.4]
  assign _GEN_0 = ~RW0_wmode;
  assign _GEN_1 = ~RW0_wmode;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {2{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    ram[initvar] = _RAND_0[43:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge RW0_clk) begin
    if(ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data; // @[:anonymous source@1266.4]
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & _GEN_0;
    if (RW0_en & _GEN_0) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
endmodule
